`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ECE-Illinois
// Engineer: Zuofu Cheng
// 
// Create Date: 06/08/2023 12:21:05 PM
// Design Name: 
// Module Name: hdmi_text_controller_v1_0_AXI
// Project Name: ECE 385 - hdmi_text_controller
// Target Devices: 
// Tool Versions: 
// Description: 
// This is a modified version of the Vivado template for an AXI4-Lite peripheral,
// rewritten into SystemVerilog for use with ECE 385.
// 
// Dependencies: 
// 
// Revision:
// Revision 0.02 - File modified to be more consistent with generated template
// Revision 11/18 - Made comments less confusing
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


`timescale 1 ns / 1 ps

module hdmi_text_controller_v1_0_AXI #
(

    // Parameters of Axi Slave Bus Interface S_AXI
    // Modify parameters as necessary for access of full VRAM range

    // Width of S_AXI data bus
    parameter integer C_S_AXI_DATA_WIDTH	= 32,
    // Width of S_AXI address bus
    parameter integer C_S_AXI_ADDR_WIDTH	= 16
)
(
    // Users to add ports here

//    output logic [31:0] controlData,
    input logic [C_S_AXI_ADDR_WIDTH-1 : 0] calcAddr,
    output logic [31:0] calcData,

   input logic [3:0] FGD_idx,
   input logic [3:0] BGD_idx,                         //used in Lab 7.2
   output logic [11:0] FGD_color,
   output logic [11:0] BGD_color,

    // User ports ends

    // Global Clock Signal
    input logic  S_AXI_ACLK,
    // Global Reset Signal. This Signal is Active LOW
    input logic  S_AXI_ARESETN,
    // Write address (issued by master, acceped by Slave)
    input logic [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
    // Write channel Protection type. This signal indicates the
        // privilege and security level of the transaction, and whether
        // the transaction is a data access or an instruction access.
    input logic [2 : 0] S_AXI_AWPROT,
    // Write address valid. This signal indicates that the master signaling
        // valid write address and control information.
    input logic  S_AXI_AWVALID,
    // Write address ready. This signal indicates that the slave is ready
        // to accept an address and associated control signals.
    output logic  S_AXI_AWREADY,
    // Write data (issued by master, acceped by Slave) 
    input logic [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_WDATA,
    // Write strobes. This signal indicates which byte lanes hold
        // valid data. There is one write strobe bit for each eight
        // bits of the write data bus.    
    input logic [(C_S_AXI_DATA_WIDTH/8)-1 : 0] S_AXI_WSTRB,
    // Write valid. This signal indicates that valid write
        // data and strobes are available.
    input logic  S_AXI_WVALID,
    // Write ready. This signal indicates that the slave
        // can accept the write data.
    output logic  S_AXI_WREADY,
    // Write response. This signal indicates the status
        // of the write transaction.
    output logic [1 : 0] S_AXI_BRESP,
    // Write response valid. This signal indicates that the channel
        // is signaling a valid write response.
    output logic  S_AXI_BVALID,
    // Response ready. This signal indicates that the master
        // can accept a write response.
    input logic  S_AXI_BREADY,
    // Read address (issued by master, acceped by Slave)
    input logic [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
    // Protection type. This signal indicates the privilege
        // and security level of the transaction, and whether the
        // transaction is a data access or an instruction access.
    input logic [2 : 0] S_AXI_ARPROT,
    // Read address valid. This signal indicates that the channel
        // is signaling valid read address and control information.
    input logic  S_AXI_ARVALID,
    // Read address ready. This signal indicates that the slave is
        // ready to accept an address and associated control signals.
    output logic  S_AXI_ARREADY,
    // Read data (issued by slave)
    output logic [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_RDATA,
    // Read response. This signal indicates the status of the
        // read transfer.
    output logic [1 : 0] S_AXI_RRESP,
    // Read valid. This signal indicates that the channel is
        // signaling the required read data.
    output logic  S_AXI_RVALID,
    // Read ready. This signal indicates that the master can
        // accept the read data and response information.
    input logic  S_AXI_RREADY
);

// AXI4LITE signals
logic  [C_S_AXI_ADDR_WIDTH-1 : 0] 	axi_awaddr;
logic  axi_awready;
logic  axi_wready;
logic  [1 : 0] 	axi_bresp;
logic  axi_bvalid;
logic  [C_S_AXI_ADDR_WIDTH-1 : 0] 	axi_araddr;
logic  axi_arready;
logic  [C_S_AXI_DATA_WIDTH-1 : 0] 	axi_rdata;
logic  [1 : 0] 	axi_rresp;
logic  	axi_rvalid;

// Example-specific design signals
// local parameter for addressing 32 bit / 64 bit C_S_AXI_DATA_WIDTH
// ADDR_LSB is used for addressing 32/64 bit registers/memories
// ADDR_LSB = 2 for 32 bits (n downto 2)
// ADDR_LSB = 3 for 64 bits (n downto 3)
localparam integer ADDR_LSB = (C_S_AXI_DATA_WIDTH/32) + 1;
localparam integer OPT_MEM_ADDR_BITS = 9;
//----------------------------------------------
//-- Signals for user logic register space example
//------------------------------------------------
//-- Number of Slave Registers 4
//logic [C_S_AXI_DATA_WIDTH-1:0]	slv_reg0;
//logic [C_S_AXI_DATA_WIDTH-1:0]	slv_reg1;
//logic [C_S_AXI_DATA_WIDTH-1:0]	slv_reg2;
//logic [C_S_AXI_DATA_WIDTH-1:0]	slv_reg3;
//
//Note: the provided Verilog template had the registered declared as above, but in order to give 
//students a hint we have replaced the 4 individual registers with an unpacked array of packed logic. 
//Note that you as the student will still need to extend this to the full register set needed for the lab.
//logic [C_S_AXI_DATA_WIDTH-1:0] slv_regs[601];
logic	 slv_reg_rden;
logic	 slv_reg_wren;
logic [C_S_AXI_DATA_WIDTH-1:0]	 reg_data_out;
//integer	 byte_index;
logic	 aw_en;

// I/O Connections assignments

assign S_AXI_AWREADY	= axi_awready;
assign S_AXI_WREADY	= axi_wready;
assign S_AXI_BRESP	= axi_bresp;
assign S_AXI_BVALID	= axi_bvalid;
assign S_AXI_ARREADY = axi_arready;
assign S_AXI_RDATA	= axi_rdata;
assign S_AXI_RRESP	= axi_rresp;
assign S_AXI_RVALID	= axi_rvalid;

// BRAM Connections
localparam integer BRAM_ADDR_WIDTH = 11;

logic [BRAM_ADDR_WIDTH-1:0] addra, addrb;
logic [C_S_AXI_DATA_WIDTH-1:0] dina, douta, doutb;
logic [3:0] wea;
logic ena, ena_wr, ena_rd;
//assign ena = ena_wr | ena_rd;
assign ena = slv_reg_wren | slv_reg_rden;

logic [10:0] tempAddr;
assign tempAddr = calcAddr;
assign addrb = calcAddr;
assign calcData = doutb;
//assign controlData = 32'h001F6000;  //hard coded for lab 7.1 (not needed for lab 7.2)

//Lab 7.2 stuff
logic [C_S_AXI_DATA_WIDTH-1:0] palette[16];
logic [11:0] Fcolor, Bcolor;
assign FGD_color = Fcolor;
assign BGD_color = Bcolor;

always_comb
begin
   Fcolor = palette[FGD_idx][11:0];
   Bcolor = palette[BGD_idx][11:0];
end



//BRAM instantiation

blk_mem_gen_0 memory (
        .addra(addra),                                          //addres to be writen to or read from
        .clka(S_AXI_ACLK),                                      //clock for synchornization
        .dina(dina),                                            //data to write into memory
        .ena(ena),       //ena_wr | ena_rd                      //enable port (must be high for both read and write operations)
        .wea(wea),                                              //Write_enable (which bytes of din do we want to write to memory, the STRB signal)
        .douta(douta),                                          //data read from memory
        
        .addrb(addrb),          //addrb, comes from calculating what grid spot we are displaying so need to get the data for that space
        .clkb(S_AXI_ACLK),
        .dinb(32'h00000000),    //never write to memory so always 0's
        .enb(1'b1),             //always reading so can just put 1
        .web(4'b0000),          //always read so has to be 4'b0000
        .doutb(doutb)           //contains 2 "spaces", Inversion bit, 7 bits of glyph data, 4 bits of FGD color index, 4 bits of BGD color index
);

always_ff @(posedge S_AXI_ACLK)
begin
    dina <= S_AXI_WDATA;
end

//hardcode palette registers
//always_comb
//begin
//    palette[0] = 12'h000;
//    palette[1] = 12'h00F;
//    palette[2] = 12'h0F0;
//    palette[3] = 12'h0FF;
//    palette[4] = 12'hF00;
//    palette[5] = 12'hF0F;
//    palette[6] = 12'hFF0;
//    palette[7] = 12'hFFF;
//    palette[8] = 12'h007;
//    palette[9] = 12'h070;
//    palette[10] = 12'h077;
//    palette[11] = 12'h700;
//    palette[12] = 12'h707;
//    palette[13] = 12'h770;
//    palette[14] = 12'h777;
//    palette[15] = 12'h333;
//    palette[16] = 12'hBBB;
//end



// Implement axi_awready generation
// axi_awready is asserted for one S_AXI_ACLK clock cycle when both
// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_awready is
// de-asserted when reset is low.

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_awready <= 1'b0;
      aw_en <= 1'b1;
    end 
  else
    begin    
      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en)
        begin
          // slave is ready to accept write address when 
          // there is a valid write address and write data
          // on the write address and data bus. This design 
          // expects no outstanding transactions. 
          axi_awready <= 1'b1;
          aw_en <= 1'b0;
        end
        else if (S_AXI_BREADY && axi_bvalid)
            begin
              aw_en <= 1'b1;
              axi_awready <= 1'b0;
            end
      else           
        begin
          axi_awready <= 1'b0;
        end
    end 
end       

// Implement axi_awaddr latching
// This process is used to latch the address when both 
// S_AXI_AWVALID and S_AXI_WVALID are valid. 

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_awaddr <= 0;
    end 
  else
    begin    
      if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en)
        begin
          // Write Address latching 
          axi_awaddr <= S_AXI_AWADDR;
        end
    end 
end       

// Implement axi_wready generation
// axi_wready is asserted for one S_AXI_ACLK clock cycle when both
// S_AXI_AWVALID and S_AXI_WVALID are asserted. axi_wready is 
// de-asserted when reset is low. 

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_wready <= 1'b0;
    end 
  else
    begin    
      if (~axi_wready && S_AXI_WVALID && S_AXI_AWVALID && aw_en )
        begin
          // slave is ready to accept write data when 
          // there is a valid write address and write data
          // on the write address and data bus. This design 
          // expects no outstanding transactions. 
          axi_wready <= 1'b1;
        end
      else
        begin
          axi_wready <= 1'b0;
        end
    end 
end       

// Implement memory mapped register select and write logic generation
// The write data is accepted and written to memory mapped registers when
// axi_awready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted. Write strobes are used to
// select byte enables of slave registers while writing.
// These registers are cleared when reset (active low) is applied.
// Slave register write enable is asserted when valid address and data are available
// and the slave is ready to accept the write address and write data.
assign slv_reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;
logic [11:0] write_addr;
logic [11:0] read_addr;
assign write_addr = S_AXI_AWADDR[2*ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB]; // 13 : 2
assign read_addr = S_AXI_ARADDR[2*ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB]; // 13 : 2

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 ) // maybe include
    begin
        palette[0] = 12'h000;   //on reset go to these random colors
        palette[1] = 12'h000;       //change to go to all 0's later
        palette[2] = 12'h000;
        palette[3] = 12'h000;
        palette[4] = 12'h000;
        palette[5] = 12'h000;
        palette[6] = 12'h000;
        palette[7] = 12'h000;
        palette[8] = 12'h000;
        palette[9] = 12'h000;
        palette[10] = 12'h000;
        palette[11] = 12'h000;
        palette[12] = 12'h000;
        palette[13] = 12'h000;
        palette[14] = 12'h000;
        palette[15] = 12'h000;
        palette[16] = 12'h000;
      //  axi_rdata <= 32'h00000000;
      //  for (integer i = 0; i < 1200; i++)
      //  begin
      //     addra <= i;                //set address (loops thru all 1200 memory addresses)
      //     wea <= 4'b1111;            //write all 4 bytes
      //     dina <= 32'h00000000;      //set to 0's
      //  end
    end
  else begin
    if (slv_reg_wren)
      begin
        if(S_AXI_AWADDR[13]) // change ot 13
          begin
           palette[write_addr[3:0]] <= S_AXI_WDATA;       //lab 7.2 stuff
          end
//        addra <= axi_awaddr[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB];
//        wea <= S_AXI_WSTRB;
//        dina <= S_AXI_WDATA;

////        for ( byte_index = 0; byte_index <= (C_S_AXI_DATA_WIDTH/8)-1; byte_index = byte_index+1 )
////         if ( S_AXI_WSTRB[byte_index] == 1 ) begin
////            // Respective byte enables are asserted as per write strobes, note the use of the index part select operator
////            // '+:', you will need to understand how this operator works.
////            slv_regs[axi_awaddr[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB]][(byte_index*8) +: 8] <= S_AXI_WDATA[(byte_index*8) +: 8];
////          end  
      end
//    else if (slv_reg_rden)
//        begin
//          addra <= axi_araddr[ADDR_LSB+OPT_MEM_ADDR_BITS:ADDR_LSB];
//          wea <= 4'b0000;
//          ena_rd <= 1'b1;
////          axi_rdata <= reg_data_out;     // register read data
//        end
  end
end

//always_ff @(posedge S_AXI_ACLK)
//begin
//    delay <= 1'b0;
//    if(ena_rd)
//    begin
//        delay <= 1'b1;
//    end
//end

//logic delay;
//always_ff @(posedge S_AXI_ACLK)
//begin
//    if(delay)
//    begin
//        axi_rdata <= reg_data_out;
//    end
//end

// Implement write response logic generation
// The write response and response valid signals are asserted by the slave 
// when axi_wready, S_AXI_WVALID, axi_wready and S_AXI_WVALID are asserted.  
// This marks the acceptance of address and indicates the status of 
// write transaction.

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_bvalid  <= 0;
      axi_bresp   <= 2'b0;
    end 
  else
    begin    
      if (axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID)
        begin
          // indicates a valid write response is available
          axi_bvalid <= 1'b1;
          axi_bresp  <= 2'b0; // 'OKAY' response 
        end                   // work error responses in future
      else
        begin
          if (S_AXI_BREADY && axi_bvalid) 
            //check if bready is asserted while bvalid is high) 
            //(there is a possibility that bready is always asserted high)   
            begin
              axi_bvalid <= 1'b0; 
            end  
        end
    end
end   

// Implement axi_arready generation
// axi_arready is asserted for one S_AXI_ACLK clock cycle when
// S_AXI_ARVALID is asserted. axi_awready is 
// de-asserted when reset (active low) is asserted. 
// The read address is also latched when S_AXI_ARVALID is 
// asserted. axi_araddr is reset to zero on reset assertion.

always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_arready <= 1'b0;
      axi_araddr  <= 32'b0;
    end 
  else
    begin    
      if (~axi_arready && S_AXI_ARVALID)
        begin
          // indicates that the slave has acceped the valid read address
          axi_arready <= 1'b1;
          // Read address latching
          axi_araddr  <= S_AXI_ARADDR;
        end
      else
        begin
          axi_arready <= 1'b0;
        end
    end 
end       

// Implement axi_arvalid generation
// axi_rvalid is asserted for one S_AXI_ACLK clock cycle when both 
// S_AXI_ARVALID and axi_arready are asserted. The slave registers 
// data are available on the axi_rdata bus at this instance. The 
// assertion of axi_rvalid marks the validity of read data on the 
// bus and axi_rresp indicates the status of read transaction.axi_rvalid 
// is deasserted on reset (active low). axi_rresp and axi_rdata are 
// cleared to zero on reset (active low).  
logic delay;
always_ff @(posedge S_AXI_ACLK)
begin
    delay <= 1'b0;
    if(slv_reg_rden)
    begin
        delay <= 1'b1;
    end
end


always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_rvalid <= 0;
      axi_rresp  <= 0;
    end 
  else
    begin    
      if (delay) //(axi_arready && S_AXI_ARVALID && ~axi_rvalid)
        begin
          // Valid read data is available at the read data bus
          axi_rvalid <= 1'b1;
          axi_rresp  <= 2'b0; // 'OKAY' response
        end   
      else if (axi_rvalid && S_AXI_RREADY)
        begin
          // Read data is accepted by the master
          axi_rvalid <= 1'b0;
        end                
    end
end    

// Implement memory mapped register select and read logic generation
// Slave register read enable is asserted when valid address is available
// and the slave is ready to accept the read address.
assign slv_reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;
//always_comb
//begin
//      // Address decoding for reading registers
//     reg_data_out = douta;
//end
logic [C_S_AXI_DATA_WIDTH-1 : 0] assigned_data;
always_comb
begin
  if (S_AXI_ARADDR[13])   //(S_AXI_ARADDR[13] && read_addr[3:0] < 16)
  begin
    assigned_data <= palette[read_addr[3:0]];
  end else
  begin
    assigned_data <= douta;
  end
end
// Output register or memory read data
always_ff @( posedge S_AXI_ACLK )
begin
  if ( S_AXI_ARESETN == 1'b0 )
    begin
      axi_rdata  <= 0;
    end 
  else
    begin    
      // When there is a valid read address (S_AXI_ARVALID) with 
      // acceptance of read address by the slave (axi_arready), 
      // output the read dada 
    //  if (slv_reg_rden && S_AXI_ARADDR[13])
    //  begin
    //    axi_rdata <= palette[read_addr[3:0]];
    //  end 
      if (delay)
        begin
          axi_rdata <= assigned_data;     // register read data
        end 
    end
end    



// Add user logic here
always_comb
begin
      if(slv_reg_wren && ~S_AXI_AWADDR[13])
      begin
          addra = axi_awaddr[ADDR_LSB+1+OPT_MEM_ADDR_BITS:ADDR_LSB];
          wea = S_AXI_WSTRB;
      end
      else if (slv_reg_rden)
      begin
          addra = axi_araddr[ADDR_LSB+1+OPT_MEM_ADDR_BITS:ADDR_LSB];
          wea = 4'h0;
      end
end

// User logic ends

endmodule
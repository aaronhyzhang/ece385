`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/26/2025 09:49:51 PM
// Design Name: 
// Module Name: digit_rom
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module digit_rom (
  input  logic [3:0] digit,  // 0-9
  input  logic [3:0] row,    // 0-15
  output logic [7:0] bits    // one byte per row
);

  always_comb begin
    unique case (digit)
      // ?????????????????????????????????????????????????????????????????????????
      4'd0: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 00111100
        4'd2:  bits = 8'b01111100; // 01000010
        4'd3:  bits = 8'b11000110; // 10000001
        4'd4:  bits = 8'b11000110;
        4'd5:  bits = 8'b11001110;
        4'd6:  bits = 8'b11011110;
        4'd7:  bits = 8'b11110110;
        4'd8:  bits = 8'b11100110;
        4'd9:  bits = 8'b11000110;
        4'd10: bits = 8'b11000110;
        4'd11: bits = 8'b01111100;
        4'd12: bits = 8'b00000000;
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      4'd1: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 00001000
        4'd2:  bits = 8'b00011000; // 00011000
        4'd3:  bits = 8'b00111000; // 00101000
        4'd4:  bits = 8'b01111000;
        4'd5:  bits = 8'b00011000;
        4'd6:  bits = 8'b00011000;
        4'd7:  bits = 8'b00011000;
        4'd8:  bits = 8'b00011000;
        4'd9:  bits = 8'b00011000;
        4'd10: bits = 8'b00011000;
        4'd11: bits = 8'b01111110;
        4'd12: bits = 8'b00000000; // 00111110
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      4'd2: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 00111100
        4'd2:  bits = 8'b01111100; // 01000010
        4'd3:  bits = 8'b11000110; // 00000010
        4'd4:  bits = 8'b00000110; // 00000100
        4'd5:  bits = 8'b00001100; // 00001000
        4'd6:  bits = 8'b00011000; // 00010000
        4'd7:  bits = 8'b00110000; // 00100000
        4'd8:  bits = 8'b01100000; // 01000000
        4'd9:  bits = 8'b11000000;
        4'd10: bits = 8'b11000110; // 01000010
        4'd11: bits = 8'b11111110; // 00111110
        4'd12: bits = 8'b00000000; // 00111110
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      4'd3: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 00111100
        4'd2:  bits = 8'b01111100; // 01000010
        4'd3:  bits = 8'b11000110; // 00000010
        4'd4:  bits = 8'b00000110;
        4'd5:  bits = 8'b00000110; // 00011100
        4'd6:  bits = 8'b00111100;
        4'd7:  bits = 8'b00000110;
        4'd8:  bits = 8'b00000110;
        4'd9:  bits = 8'b00000110;
        4'd10: bits = 8'b11000110;
        4'd11: bits = 8'b01111100;
        4'd12: bits = 8'b00000000; // 00111110
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      4'd4: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 00000100
        4'd2:  bits = 8'b00001100; // 00001100
        4'd3:  bits = 8'b00011100; // 00010100
        4'd4:  bits = 8'b00111100; // 00100100
        4'd5:  bits = 8'b01101100; // 01000100
        4'd6:  bits = 8'b11001100; // 01111110
        4'd7:  bits = 8'b11111110;
        4'd8:  bits = 8'b00001100;
        4'd9:  bits = 8'b00001100;
        4'd10: bits = 8'b00001100;
        4'd11: bits = 8'b00011110; // 00001111
        4'd12: bits = 8'b00000000; // 00111110
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      4'd5: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 01111110
        4'd2:  bits = 8'b11111110; // 01100000
        4'd3:  bits = 8'b11000000;
        4'd4:  bits = 8'b11000000; // 01111100
        4'd5:  bits = 8'b11000000; // 00000110
        4'd6:  bits = 8'b11111100; // 00000010
        4'd7:  bits = 8'b00000110;
        4'd8:  bits = 8'b00000110;
        4'd9:  bits = 8'b00000110; // 01000010
        4'd10: bits = 8'b11000110;
        4'd11: bits = 8'b01111100; // 00111100
        4'd12: bits = 8'b00000000; // 00111110
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      4'd6: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 00111100
        4'd2:  bits = 8'b00111000; // 01000010
        4'd3:  bits = 8'b01100000; // 01000000
        4'd4:  bits = 8'b11000000;
        4'd5:  bits = 8'b11000000; // 01111100
        4'd6:  bits = 8'b11111100; // 01100110
        4'd7:  bits = 8'b11000110; // 01100011
        4'd8:  bits = 8'b11000110;
        4'd9:  bits = 8'b11000110;
        4'd10: bits = 8'b11000110;
        4'd11: bits = 8'b01111100; // 00111110
        4'd12: bits = 8'b00000000; // 00111110
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      4'd7: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 01111110
        4'd2:  bits = 8'b11111110; // 01000010
        4'd3:  bits = 8'b11000110; // 00000010
        4'd4:  bits = 8'b00000110; // 00000100
        4'd5:  bits = 8'b00000110;
        4'd6:  bits = 8'b00001100;
        4'd7:  bits = 8'b00011000;
        4'd8:  bits = 8'b00110000;
        4'd9:  bits = 8'b00110000;
        4'd10: bits = 8'b00110000;
        4'd11: bits = 8'b00110000;
        4'd12: bits = 8'b00000000; // 00111110
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      4'd8: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 00111100
        4'd2:  bits = 8'b01111100; // 01100110
        4'd3:  bits = 8'b11000110;
        4'd4:  bits = 8'b11000110; // 00111100
        4'd5:  bits = 8'b11000110;
        4'd6:  bits = 8'b01111100;
        4'd7:  bits = 8'b11000110;
        4'd8:  bits = 8'b11000110;
        4'd9:  bits = 8'b11000110;
        4'd10: bits = 8'b11000110;
        4'd11: bits = 8'b01111100;
        4'd12: bits = 8'b00000000; // 00111110
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      4'd9: unique case (row)
        4'd0:  bits = 8'b00000000;
        4'd1:  bits = 8'b00000000; // 00111100
        4'd2:  bits = 8'b01111100; // 01100110
        4'd3:  bits = 8'b11000110;
        4'd4:  bits = 8'b11000110;
        4'd5:  bits = 8'b11000110; // 00111110
        4'd6:  bits = 8'b01111110; // 00000110
        4'd7:  bits = 8'b00000110;
        4'd8:  bits = 8'b00000110;
        4'd9:  bits = 8'b00000110;
        4'd10: bits = 8'b00001100;
        4'd11: bits = 8'b01111000;
        4'd12: bits = 8'b00000000; // 00111110
        4'd13: bits = 8'b00000000;
        4'd14: bits = 8'b00000000;
        4'd15: bits = 8'b00000000;
        default: bits = 8'h00;
      endcase

      // ?????????????????????????????????????????????????????????????????????????
      default: bits = 8'h00;
    endcase
  end

endmodule

